module tb_SingleCPU;
reg [31:0] Addr_in;
reg clk;
wire [31:0] Addr_o;
// wire [31:0]alu_result;
// wire ALUSrc;
// wire [31:0]mux32b1_out;
// wire [31:0]dm_out;
integer i;

SingleCPU uut(
    Addr_in,
    clk,
    Addr_o
    // alu_result,
    // ALUSrc
    // mux32b1_out,
    // dm_out
);

initial begin
    i <= 0;
    clk <= 0;
    #10
    clk <= !clk;
    for(i=0;i<64;i=i+4)begin
        #10
        clk <= !clk;
        #10
        clk <= !clk;
        Addr_in <= i;
    end


end


endmodule